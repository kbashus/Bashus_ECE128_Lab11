`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 11/27/2023 04:58:16 PM
// Design Name: 
// Module Name: RegisterNbit
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module RegisterNbit(D, Q,  L, R, clock);

    parameter N = 4; // number of bits

    output reg [N-1:0]Q; // registered output
    input [N-1:0]D; // data input
    input L; // load enable
    input R; // positive logic asynchronous reset
    input clock; // positive edge clock
    
                 
    always @(posedge clock or posedge R) begin

    if(R)
        Q <= 0;
    else if(L)
        Q <= D;
    else
        Q <= Q;
end

endmodule
